library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity temp is
	port(
			DQ		    :inout STD_LOGIC;  					 -- DS18B20??????
			inclk       :in std_logic;						 --??????
			current_temp:out std_logic_vector(10 downto 0)   --?????????4?????????7??????
		);
end entity;

architecture Behavior of temp is

	--????????0xcc??????????????0xcc
	constant cmd_0xcc_0x44:std_logic_vector(15 downto 0):="00110011"&"00100010";   --ROM???~0xcc ?0x44
	constant cmd_0xcc_0xbe:std_logic_vector(15 downto 0):="00110011"&"01111101";   --ROM???~0xcc ?0xbe
	signal temp1,temp2:std_logic_vector(7 downto 0);    --???????
	signal nflag:std_logic;    --????????????????????	
	signal clk:std_logic;   --??????????	
	signal count:std_logic_vector(4 downto 0); --???????
	--???????	
	begin
		process(inclk)
		begin
			if rising_edge(inclk) then	
				if (count="11010") then --1MHZ
					clk<=not clk;
					count<="00000";
				else
					count<=count+1;
				end if;
			end if;
		end process;

	process(clk)
		variable count1:std_logic_vector(10 downto 0);   --???1???DS18B20????????????
		variable count2:std_logic_vector(9 downto 0);   --???2????DS18B20????????????
		variable count3:std_logic_vector(7 downto 0);   --???3????DS18B20????????????

		variable i:integer range -1 to 15:=15;   --???????
		variable init:integer range 0 to 1:=0;   --???????
		variable j:integer range 0 to 8:=0;      --??????????
		variable k:integer range 0 to 1:=0;      --???????????
		variable state:integer range 0 to 2:=0;   --?????0????1,1????2,2?????

		variable temp:std_logic_vector(7 downto 0);
		begin
			if rising_edge(clk) then
				if state=0 then
					if init=1 then   --????????????
						count2:=count2+1;
					if count2="0000000001" then   --?????
						DQ<='0';
					elsif count2="0000001100" then   --?15us??????????
						DQ<=cmd_0xcc_0x44(i);
					elsif count2="0001011010" then   --?????15us~60us??DS18B20?????????90us
						DQ<='1';
					elsif count2="1010110100" then   --???1us???????????????
						count2:="0000000000";   --?????
						i:=i-1;   --??1????
						if i=-1 then    --??????????????????????????????????1??????2
							i:=15;init:=0;state:=1;
						end if;
					end if;
				else   --init=0??????
					count1:=count1+1;
					if count1="000000000001" then
						DQ<='1';
					elsif count1="000000000011" then   --??
						DQ<='0';
					elsif count1="01010111100" then   --??????????????480us????500us
						DQ<='1';
					elsif count1="01011011010" then   --??15us~60us???????30us?530??????????DS18B20??????
						DQ<='Z';
					elsif count1="01111001010" then   --?????60us~240us?830????
						DQ<='1';
					elsif count1="10000000000" then   --??????960us????1024us
						init:=1;
						count1:="00000000000";   --???????????????????1????????????????
					end if;
				end if;
			elsif (state=1) then   --state=1????2
				if init=1 then
					count2:=count2+1;
					if count2="0000000001" then
						DQ<='0';
					elsif count2="0000001100" then
						DQ<=cmd_0xcc_0xbe(i);
					elsif count2="0001011010" then
						DQ<='1';
					elsif count2="0001011100" then
						count2:="0000000000";
						i:=i-1;
						if i=-1 then
							i:=15;
							init:=0;
							state:=2;
						end if;
					end if;
				else
					count1:=count1+1;
					if count1="000000000001" then
						DQ<='1';
					elsif count1="000000000011" then   --??
						DQ<='0';
					elsif count1="01010111100" then   --??????????????480us????500us
						DQ<='1';
					elsif count1="01011011010" then   --??15us~60us???????30us?530??????????DS18B20??????
						DQ<='Z';
					elsif count1="01111001010" then   --?????60us~240us?830????
						DQ<='1';
					elsif count1="10000000000" then   --??????960us????1024us
						init:=1;
						count1:="00000000000";   --???????????????????1????????????????
					end if;
				end if;
			else    --state=2?????
				if k=0 then   --k=0??????????????
					count3:=count3+1;
					if count3="00000001" then
						DQ<='0';
					elsif count3="00000100" then   --?????1us??????
						DQ<='Z';
					elsif count3="00001101" then   --???15us?????
						temp(j):=DQ;
					elsif count3="01010000" then   --?????60us????80us
						DQ<='1';
					elsif count3="01010010" then   --?????
						count3:="00000000";
						j:=j+1;   --??????
						if j=8 then   --???
							j:=0;   --?0
							k:=1;   --??2??
							temp1<=temp;
						end if;
					end if;
				else   --k=1 ??2??
					count3:=count3+1;
						if count3="00000001" then
							DQ<='0';
						elsif count3="00000100" then
							DQ<='Z';
						elsif count3="00001101" then
							temp(j):=DQ;
						elsif count3="01010000" then
							DQ<='1';
						elsif count3="01010010" then
							count3:="00000000";
							j:=j+1;
							if j=8 then
								j:=0;
								k:=0;
								state:=0;   --??????????????
								if (temp and "11111000")="11111000" then   --?????????????
									temp:=(not temp);
									temp1<=(not temp1)+1;
								if temp1="0000000" then 
									temp:=temp+1;
								end if;
									nflag<='1';   --?????
								else
									nflag<='0';
								end if;
							current_temp<=temp(2 downto 0) & temp1;   --????temp_value2??5??temp_value1
							end if;
						end if;
					end if;
				end if;
			end if;
		end process;
end  Behavior;

